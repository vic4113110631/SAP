/*
su    Fun
00   +
01   -
10   AND
11   OR
*/
module ALU( ALU_Out, A_in, B_in, su, eu);
 output ALU_Out;
 input A_in, B_in, su, eu;
 
 wire [7:0] ALU_Out;
 wire [7:0] A_in, B_in;
 wire [1:0] su;
 wire	    eu;
 
 reg       CarryOut;
 reg [6:0] Sum;
 
 always@(A_in or B_in or su)
 begin
   case(su)
     2'b00: {CarryOut, Sum} <= A_in + B_in;
     2'b01: {CarryOut, Sum} <= A_in - B_in;
     2'b10: {CarryOut, Sum} <= A_in & B_in;
     2'b11: {CarryOut, Sum} <= A_in | B_in;
   endcase
 end

 assign ALU_Out = eu ? {CarryOut, Sum} : 8'bz;

endmodule
